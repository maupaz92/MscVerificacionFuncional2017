class estimulo3;

endclass