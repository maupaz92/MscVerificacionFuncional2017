


program test(
	interface driver_port,
	interface monitor_port,
	interface config_port
);


	environment test_bench_environment;













endprogram











