


program test(
	interface driver_port,
	interface monitor_port,
	interface config_port
);


	environment test_bench_environment;
	
	initial begin
		
		test_bench_environment = new();
	
	end 













endprogram











