class estimulo2;

endclass